module uart_top(
    input clk, // The master clock for this module
    input rst_n, // Synchronous reset.
    input rx, // Incoming serial line
    output tx, // Outgoing serial line
    output [7:0] rx_byte, // Byte received
	 output debug_output
);

//uart
logic is_receiving;
logic is_transmitting;
logic recv_error;
logic received;
logic transmit;
logic [7:0] tx_byte;

logic received_q, received_d;
logic [7:0] rx_byte_internal;
logic [7:0] rx_store_q, rx_store_d;

//debug
logic [7:0]	debug_q,debug_d;

  always_comb begin
    rx_store_d = rx_store_q;
	 received_d = received;
	 debug_d 	= debug_q;
    if ( received ) begin
	  rx_store_d = rx_byte_internal;
	  debug_d 	 = !debug_q;
    end
  end 

  always_ff @ (posedge clk or negedge rst_n) begin
    if (!rst_n) begin
	    rx_store_q <=	'0; 
		 received_q <= '0;
		 debug_q 	<= '0;
    end
    else begin
	    rx_store_q <= rx_store_d;
		 received_q <=	received_d;
		 debug_q 	<=	debug_d;
    end
  end
	
    uart i_uart(
        .clk(clk),
        .rst(rst_n),
        .rx(rx),
        .tx(tx),
        .transmit(received_q),
        .tx_byte(rx_store_q),
        .received(received),
        .rx_byte(rx_byte_internal),
        .is_receiving(is_receiving),
        .is_transmitting(is_transmitting),
        .recv_error(recv_error)
    );
	 
	 //assign received 		= received_q;
	 assign rx_byte 		= rx_store_q;
	 assign debug_output = debug_q;
	 
endmodule
